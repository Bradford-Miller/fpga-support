-- ------------------------------------------------
--                                               --
-- Temporary "library" to develop pad code       --
--                                               --
-- Time-stamp: <2022-05-02 14:04:44 gorbag>      --
--                                               --
-- ------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package padpkg is

end package padpkg;

package body padpkg is

end package body padpkg;
