work/regpkg.vhdl